library ieee;
use ieee.std_logic_1164.all;

package config is

  -- input file path :
  constant input_path : string :="C:\Users\Ryuuk\Desktop\Nouveau dossier\pgm\horz.pgm";
  -- output file path :
  constant output_path : string :="C:\Users\Ryuuk\Desktop\Nouveau dossier\pgm\test.pgm";
  -- image width
  constant image_width : integer := 20;

end config;
